// When this is defined, the types of TRegFile will be defined in OptimisedCompile and imported.
`define HCHAL_OPTIMISED_COMPILE
